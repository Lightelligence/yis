// Copyright (c) 2020 Lightelligence
// Description: FIFO Wrappers Interface generated from test_fifo_a.yis by YIS
