// Copyright (c) 2020 Lightelligence
// Description: Memory Wrappers Interface generated from test_mem_a.yis by YIS


///////////////////////////////////////////////////////////////////////////////
// name: rx_fifo
// doc_summary: Receive FIFO Memory
/* doc_verbose: Boring info about memories. And now
I'm on a new line
 */
// width: test_pkg_a::TRIPLE_NESTED_PARAM.value  ==>  2
// depth: 512  ==>  512
// ecc: True
// parity: False
// sram_type: 2p

module rx_fifo_mem_wrapper
(
// FIXME ports
);

// FIXME module body

endmodule : rx_fifo_mem_wrapper

///////////////////////////////////////////////////////////////////////////////
// name: tx_fifo
// doc_summary: Transimit FIFO Memory

// width: test_pkg_a::hero_write__st.width  ==>  46
// depth: 1024  ==>  1024
// ecc: False
// parity: True
// sram_type: 1p

module tx_fifo_mem_wrapper
(
// FIXME ports
);

// FIXME module body

endmodule : tx_fifo_mem_wrapper
